module cm ( 
	a,
	b,
	ma,
	me,
	i
	) ;

input [3:0] a;
input [3:0] b;
inout  ma;
inout  me;
inout  i;
