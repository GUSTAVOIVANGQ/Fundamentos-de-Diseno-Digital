module su ( 
	a,
	b,
	ci,
	s,
	cf
	) ;

input [3:0] a;
input [3:0] b;
input  ci;
inout [3:0] s;
inout  cf;
