LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY MUX IS port(
A,B : IN STD_LOGIC;
S:IN STD_LOGIC_VECTOR(2 DOWNTO 0);
Z: OUT STD_LOGIC
);
END ENTITY;

ARCHITECTURE A_MUX OF MUX IS
BEGIN
process(S)
BEGIN
CASE S IS
WHEN "000"=> Z <= A OR B;
WHEN "001"=> Z <= A AND B;
WHEN "010"=> Z <= A NOR B;
WHEN "011"=> Z <= A NAND B;
WHEN "100"=> Z <= A XOR B;
WHEN "101"=> Z <= A XNOR B;
WHEN "110"=> Z <= NOT A;
WHEN OTHERS=> Z <= NOT B;
END CASE;
END PROCESS;
END A_MUX;

