LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
ENTITY CM IS
    PORT (
        A, B : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
        MA, ME, I : OUT STD_LOGIC
    );
END ENTITY;

ARCHITECTURE A_CM OF CM IS
BEGIN
    PROCESO_COMPARACION: PROCESS (A, B)
	BEGIN
	MA<='0';
	ME<='0';
	I<='0';
	IF (A = B) THEN
	I <= '1';
	ELSIF (A > B) THEN
	MA <= '1';
	ELSE
	ME<='1';
        END IF;
    END PROCESS PROCESO_COMPARACION;
END A_CM;