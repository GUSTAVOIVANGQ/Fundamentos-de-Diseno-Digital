module su ( 
	a,
	b,
	ca,
	ci,
	di,
	s,
	do,
	cf
	) ;

input [3:0] a;
input [3:0] b;
input  ca;
input  ci;
input  di;
inout [3:0] s;
inout  do;
inout  cf;
